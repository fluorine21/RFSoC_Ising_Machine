


package rfsoc_config;

parameter gpio_w_clk_bit = 24;
parameter gpio_addr_start = 15;
parameter gpio_addr_end = 0;
parameter gpio_data_start = 16;
parameter gpio_data_end = 23;



endpackage