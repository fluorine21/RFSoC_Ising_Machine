

//Allows CPU to readback A and C fifos along with status stuff over gpio

module gpio_reader
(
	input wire clk, rst,
	
	input wire [31:0] gpio_in,
	
	output reg [15:0] gpio_out,

	
);







endmodule