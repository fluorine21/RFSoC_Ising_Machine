


module experiment_fsm(
	input wire clk, rst,
	
	//Instruction bus
	input  wire instr_axis_tdata,
	input  wire instr_axis_tvalid,
	output wire instr_axis_tready,
	
	
	
	
);




endmodule