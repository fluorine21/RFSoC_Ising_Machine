import ising_config::*;


module dl_tb();

reg clk, rst;
reg [31:0] gpio_in;

reg [255:0] adc_data_in;

reg lock_sig_active, trig_lock;

wire lock_done;
wire [15:0] setpt_out_ext//Setpoint


//scale factor
real dl_to_mzi_scale_fac = 0.01;
real mzi_to_dl_scale_fac = 100;
reg [15:0] mzi_res;
real setpt_cast;

dl
#(parameter base_addr = 0) dut
(
	clk, rst, 
	gpio_in,
	
	//Incomming ADC data
	adc_data_in,
	
	lock_sig_active,//if 1, a calibration pulse is currently being read back and must be locked to
	trig_lock,//if 1, we're actively running the fsm and trying to lock
	lock_done,//If 1, this module is not in the process of locking
	
	setpt_out_ext//Setpoint output of the lockbox
);

reg [63:0] step_num;


initial begin

	test_mzi_sim();
	
	clk <= 0;
	rst <= 1;
	gpio_in <= 0;
	adc_data_in <= 0;
	lock_sig_active <= 0;
	trig_lock <= 0;
	
	repeat(10) clk_cycle();
	rst <= 0;
	repeat(10) clk_cycle();
	rst <= 1;
	repeat(10) clk_cycle();
	
	
	//Write the max_pos_tol
	gpio_write(0,0);
	//write setpt_in;
	gpio_write(1, 1000);
	//write the initial expected value exp_val_in
	gpio_write(2, 500);
	//write the tolerance
	gpio_write(3, 10);
	//write the number of averages to take 
	gpio_write(4, 2);//this is 4 averages
	gpio_write(5, 2);//lock signal pos
	
	repeat(10) clk_cycle();
	trig_lock <= 1;
	lock_sig_active <= 1;
	
	repeat (100000) step_dl_sim();
	
end





task step_dl_sim();
begin

	//Evaluate the current MZI result and feed it into the buffer
	setpt_cast = real'(setpt_out_ext*dl_to_mzi_scale_fac);
	mzi_res = 16'(run_mzi_sim(setpt_cast, get_noise())*mzi_to_dl_scale_fac);
	//Update the ADC register going into dl
	adc_data_in <= { {1{16'h0}}, 
	// cycle the clock
	clk_cycle();

end
endtask



task get_noise(output real phase);
begin
	phase = 0;
	step_num <= step_num + 1;
end
endtask






function void test_mzi_sim();

	//$display("Running MZI test");
	automatic int outfile = $fopen("mzi_test_results.csv", "w");
	real p, res, p_max;
	p_max = 20*2*pi;
	$fwrite(outfile, "p, res\n");
	
	for(p = -1*p_max; p < p_max; p = p + 0.01) begin
		res = run_mzi_sim(p, 0);
		$fwrite(outfile, "%f, %f\n", p, res);
	end
	$display("MZI test finished!");
	$fclose(outfile);
	

endfunction





function real run_mzi_sim(input real phase1, phase2);

	automatic cmp_num E0, E1, E2, E3, E4, E5;
	automatic real sf, r_fac;

	//Define the starting electric field
	E0 = '{1,0};
	
	//first beamsplitter
	E1 = cmp_mul(E0, '{1/$sqrt(2), 0});
	E2 = cmp_mul(E0, '{0, 1/$sqrt(2)});
	
	//Phase propagation
	E3 = cmp_mul(E1, cmp_exp('{0,phase1}));
	E4 = cmp_mul(E2, cmp_exp('{0,phase2}));
	
	//Second beamsplitter first output
	E5 = cmp_add(cmp_mul(E3, '{1/$sqrt(2), 0}), cmp_mul(E4, '{0, 1/$sqrt(2)}));
	
	//multiply final output intensity by exp(|x|^2) rolloff
	sf = -1/(2*pi*10);//10 wavelengths or so
	r_fac = abs(phase1-phase2)*abs(phase1-phase2)*sf;
	
	return cmp_sqr_mag(cmp_mul(E5, cmp_exp('{r_fac, 0})));

endfunction



task clk_cycle();
begin
	#1
	clk <= 1;
	#1
	#1
	clk <= 0;
	#1
	clk <= 0;
end
endtask

task gpio_write;
input [15:0] addr;
input [7:0] data;
begin
	
	clk_cycle();
	gpio_addr <= addr;
	gpio_data <= data;
	clk_cycle();
	w_clk <= 1;
	repeat(2) clk_cycle();
	w_clk <= 0;
	repeat(5) clk_cycle();
	
end
endtask

endmodule